// System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module System (
		inout  wire       aud_vid_SDAT,       //     aud_vid.SDAT
		output wire       aud_vid_SCLK,       //            .SCLK
		input  wire       clk_clk,            //         clk.clk
		input  wire       key_0_export,       //       key_0.export
		input  wire       key_1_export,       //       key_1.export
		input  wire       key_2_export,       //       key_2.export
		input  wire       key_3_export,       //       key_3.export
		output wire [9:0] red_leds_export,    //    red_leds.export
		input  wire       reset_reset_n,      //       reset.reset_n
		output wire [6:0] seven_seg_0_export, // seven_seg_0.export
		output wire [6:0] seven_seg_1_export, // seven_seg_1.export
		output wire [6:0] seven_seg_2_export, // seven_seg_2.export
		output wire [6:0] seven_seg_3_export, // seven_seg_3.export
		output wire [6:0] seven_seg_4_export, // seven_seg_4.export
		output wire [6:0] seven_seg_5_export, // seven_seg_5.export
		input  wire [9:0] switches_export     //    switches.export
	);

	wire  [31:0] niosii_data_master_readdata;                                      // mm_interconnect_0:NIOSII_data_master_readdata -> NIOSII:d_readdata
	wire         niosii_data_master_waitrequest;                                   // mm_interconnect_0:NIOSII_data_master_waitrequest -> NIOSII:d_waitrequest
	wire         niosii_data_master_debugaccess;                                   // NIOSII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOSII_data_master_debugaccess
	wire  [18:0] niosii_data_master_address;                                       // NIOSII:d_address -> mm_interconnect_0:NIOSII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                                    // NIOSII:d_byteenable -> mm_interconnect_0:NIOSII_data_master_byteenable
	wire         niosii_data_master_read;                                          // NIOSII:d_read -> mm_interconnect_0:NIOSII_data_master_read
	wire         niosii_data_master_readdatavalid;                                 // mm_interconnect_0:NIOSII_data_master_readdatavalid -> NIOSII:d_readdatavalid
	wire         niosii_data_master_write;                                         // NIOSII:d_write -> mm_interconnect_0:NIOSII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                                     // NIOSII:d_writedata -> mm_interconnect_0:NIOSII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                               // mm_interconnect_0:NIOSII_instruction_master_readdata -> NIOSII:i_readdata
	wire         niosii_instruction_master_waitrequest;                            // mm_interconnect_0:NIOSII_instruction_master_waitrequest -> NIOSII:i_waitrequest
	wire  [18:0] niosii_instruction_master_address;                                // NIOSII:i_address -> mm_interconnect_0:NIOSII_instruction_master_address
	wire         niosii_instruction_master_read;                                   // NIOSII:i_read -> mm_interconnect_0:NIOSII_instruction_master_read
	wire         niosii_instruction_master_readdatavalid;                          // mm_interconnect_0:NIOSII_instruction_master_readdatavalid -> NIOSII:i_readdatavalid
	wire  [31:0] mm_interconnect_0_audio_video_avalon_av_config_slave_readdata;    // Audio_Video:readdata -> mm_interconnect_0:Audio_Video_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_video_avalon_av_config_slave_waitrequest; // Audio_Video:waitrequest -> mm_interconnect_0:Audio_Video_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_video_avalon_av_config_slave_address;     // mm_interconnect_0:Audio_Video_avalon_av_config_slave_address -> Audio_Video:address
	wire         mm_interconnect_0_audio_video_avalon_av_config_slave_read;        // mm_interconnect_0:Audio_Video_avalon_av_config_slave_read -> Audio_Video:read
	wire   [3:0] mm_interconnect_0_audio_video_avalon_av_config_slave_byteenable;  // mm_interconnect_0:Audio_Video_avalon_av_config_slave_byteenable -> Audio_Video:byteenable
	wire         mm_interconnect_0_audio_video_avalon_av_config_slave_write;       // mm_interconnect_0:Audio_Video_avalon_av_config_slave_write -> Audio_Video:write
	wire  [31:0] mm_interconnect_0_audio_video_avalon_av_config_slave_writedata;   // mm_interconnect_0:Audio_Video_avalon_av_config_slave_writedata -> Audio_Video:writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;              // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;             // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                 // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                    // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                   // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;               // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;                // NIOSII:debug_mem_slave_readdata -> mm_interconnect_0:NIOSII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;             // NIOSII:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOSII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;             // mm_interconnect_0:NIOSII_debug_mem_slave_debugaccess -> NIOSII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;                 // mm_interconnect_0:NIOSII_debug_mem_slave_address -> NIOSII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;                    // mm_interconnect_0:NIOSII_debug_mem_slave_read -> NIOSII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;              // mm_interconnect_0:NIOSII_debug_mem_slave_byteenable -> NIOSII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;                   // mm_interconnect_0:NIOSII_debug_mem_slave_write -> NIOSII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;               // mm_interconnect_0:NIOSII_debug_mem_slave_writedata -> NIOSII:debug_mem_slave_writedata
	wire         mm_interconnect_0_red_leds_s1_chipselect;                         // mm_interconnect_0:red_leds_s1_chipselect -> red_leds:chipselect
	wire  [31:0] mm_interconnect_0_red_leds_s1_readdata;                           // red_leds:readdata -> mm_interconnect_0:red_leds_s1_readdata
	wire   [1:0] mm_interconnect_0_red_leds_s1_address;                            // mm_interconnect_0:red_leds_s1_address -> red_leds:address
	wire         mm_interconnect_0_red_leds_s1_write;                              // mm_interconnect_0:red_leds_s1_write -> red_leds:write_n
	wire  [31:0] mm_interconnect_0_red_leds_s1_writedata;                          // mm_interconnect_0:red_leds_s1_writedata -> red_leds:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                           // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                            // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_key_0_s1_chipselect;                            // mm_interconnect_0:key_0_s1_chipselect -> key_0:chipselect
	wire  [31:0] mm_interconnect_0_key_0_s1_readdata;                              // key_0:readdata -> mm_interconnect_0:key_0_s1_readdata
	wire   [1:0] mm_interconnect_0_key_0_s1_address;                               // mm_interconnect_0:key_0_s1_address -> key_0:address
	wire         mm_interconnect_0_key_0_s1_write;                                 // mm_interconnect_0:key_0_s1_write -> key_0:write_n
	wire  [31:0] mm_interconnect_0_key_0_s1_writedata;                             // mm_interconnect_0:key_0_s1_writedata -> key_0:writedata
	wire         mm_interconnect_0_seven_seg_0_s1_chipselect;                      // mm_interconnect_0:seven_seg_0_s1_chipselect -> seven_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_readdata;                        // seven_seg_0:readdata -> mm_interconnect_0:seven_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_0_s1_address;                         // mm_interconnect_0:seven_seg_0_s1_address -> seven_seg_0:address
	wire         mm_interconnect_0_seven_seg_0_s1_write;                           // mm_interconnect_0:seven_seg_0_s1_write -> seven_seg_0:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_writedata;                       // mm_interconnect_0:seven_seg_0_s1_writedata -> seven_seg_0:writedata
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                      // mm_interconnect_0:seven_seg_1_s1_chipselect -> seven_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                        // seven_seg_1:readdata -> mm_interconnect_0:seven_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                         // mm_interconnect_0:seven_seg_1_s1_address -> seven_seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                           // mm_interconnect_0:seven_seg_1_s1_write -> seven_seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                       // mm_interconnect_0:seven_seg_1_s1_writedata -> seven_seg_1:writedata
	wire         mm_interconnect_0_seven_seg_2_s1_chipselect;                      // mm_interconnect_0:seven_seg_2_s1_chipselect -> seven_seg_2:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_readdata;                        // seven_seg_2:readdata -> mm_interconnect_0:seven_seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_2_s1_address;                         // mm_interconnect_0:seven_seg_2_s1_address -> seven_seg_2:address
	wire         mm_interconnect_0_seven_seg_2_s1_write;                           // mm_interconnect_0:seven_seg_2_s1_write -> seven_seg_2:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_writedata;                       // mm_interconnect_0:seven_seg_2_s1_writedata -> seven_seg_2:writedata
	wire         mm_interconnect_0_seven_seg_3_s1_chipselect;                      // mm_interconnect_0:seven_seg_3_s1_chipselect -> seven_seg_3:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_readdata;                        // seven_seg_3:readdata -> mm_interconnect_0:seven_seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_3_s1_address;                         // mm_interconnect_0:seven_seg_3_s1_address -> seven_seg_3:address
	wire         mm_interconnect_0_seven_seg_3_s1_write;                           // mm_interconnect_0:seven_seg_3_s1_write -> seven_seg_3:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_writedata;                       // mm_interconnect_0:seven_seg_3_s1_writedata -> seven_seg_3:writedata
	wire         mm_interconnect_0_seven_seg_4_s1_chipselect;                      // mm_interconnect_0:seven_seg_4_s1_chipselect -> seven_seg_4:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_readdata;                        // seven_seg_4:readdata -> mm_interconnect_0:seven_seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_4_s1_address;                         // mm_interconnect_0:seven_seg_4_s1_address -> seven_seg_4:address
	wire         mm_interconnect_0_seven_seg_4_s1_write;                           // mm_interconnect_0:seven_seg_4_s1_write -> seven_seg_4:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_writedata;                       // mm_interconnect_0:seven_seg_4_s1_writedata -> seven_seg_4:writedata
	wire         mm_interconnect_0_seven_seg_5_s1_chipselect;                      // mm_interconnect_0:seven_seg_5_s1_chipselect -> seven_seg_5:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_readdata;                        // seven_seg_5:readdata -> mm_interconnect_0:seven_seg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_5_s1_address;                         // mm_interconnect_0:seven_seg_5_s1_address -> seven_seg_5:address
	wire         mm_interconnect_0_seven_seg_5_s1_write;                           // mm_interconnect_0:seven_seg_5_s1_write -> seven_seg_5:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_writedata;                       // mm_interconnect_0:seven_seg_5_s1_writedata -> seven_seg_5:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                            // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:chipselect
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                              // SDRAM:readdata -> mm_interconnect_0:SDRAM_s1_readdata
	wire  [14:0] mm_interconnect_0_sdram_s1_address;                               // mm_interconnect_0:SDRAM_s1_address -> SDRAM:address
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                            // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:byteenable
	wire         mm_interconnect_0_sdram_s1_write;                                 // mm_interconnect_0:SDRAM_s1_write -> SDRAM:write
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                             // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:writedata
	wire         mm_interconnect_0_sdram_s1_clken;                                 // mm_interconnect_0:SDRAM_s1_clken -> SDRAM:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                            // mm_interconnect_0:Timer_s1_chipselect -> Timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                              // Timer:readdata -> mm_interconnect_0:Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                               // mm_interconnect_0:Timer_s1_address -> Timer:address
	wire         mm_interconnect_0_timer_s1_write;                                 // mm_interconnect_0:Timer_s1_write -> Timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                             // mm_interconnect_0:Timer_s1_writedata -> Timer:writedata
	wire         mm_interconnect_0_key_1_s1_chipselect;                            // mm_interconnect_0:key_1_s1_chipselect -> key_1:chipselect
	wire  [31:0] mm_interconnect_0_key_1_s1_readdata;                              // key_1:readdata -> mm_interconnect_0:key_1_s1_readdata
	wire   [1:0] mm_interconnect_0_key_1_s1_address;                               // mm_interconnect_0:key_1_s1_address -> key_1:address
	wire         mm_interconnect_0_key_1_s1_write;                                 // mm_interconnect_0:key_1_s1_write -> key_1:write_n
	wire  [31:0] mm_interconnect_0_key_1_s1_writedata;                             // mm_interconnect_0:key_1_s1_writedata -> key_1:writedata
	wire         mm_interconnect_0_key_2_s1_chipselect;                            // mm_interconnect_0:key_2_s1_chipselect -> key_2:chipselect
	wire  [31:0] mm_interconnect_0_key_2_s1_readdata;                              // key_2:readdata -> mm_interconnect_0:key_2_s1_readdata
	wire   [1:0] mm_interconnect_0_key_2_s1_address;                               // mm_interconnect_0:key_2_s1_address -> key_2:address
	wire         mm_interconnect_0_key_2_s1_write;                                 // mm_interconnect_0:key_2_s1_write -> key_2:write_n
	wire  [31:0] mm_interconnect_0_key_2_s1_writedata;                             // mm_interconnect_0:key_2_s1_writedata -> key_2:writedata
	wire         mm_interconnect_0_key_3_s1_chipselect;                            // mm_interconnect_0:key_3_s1_chipselect -> key_3:chipselect
	wire  [31:0] mm_interconnect_0_key_3_s1_readdata;                              // key_3:readdata -> mm_interconnect_0:key_3_s1_readdata
	wire   [1:0] mm_interconnect_0_key_3_s1_address;                               // mm_interconnect_0:key_3_s1_address -> key_3:address
	wire         mm_interconnect_0_key_3_s1_write;                                 // mm_interconnect_0:key_3_s1_write -> key_3:write_n
	wire  [31:0] mm_interconnect_0_key_3_s1_writedata;                             // mm_interconnect_0:key_3_s1_writedata -> key_3:writedata
	wire         irq_mapper_receiver0_irq;                                         // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                         // key_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                         // Timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                         // key_1:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                         // key_2:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                         // key_3:irq -> irq_mapper:receiver5_irq
	wire  [31:0] niosii_irq_irq;                                                   // irq_mapper:sender_irq -> NIOSII:irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [Audio_Video:reset, NIOSII:reset_n, SDRAM:reset, Timer:reset_n, irq_mapper:reset, key_0:reset_n, key_1:reset_n, key_2:reset_n, key_3:reset_n, mm_interconnect_0:NIOSII_reset_reset_bridge_in_reset_reset, red_leds:reset_n, rst_translator:in_reset, seven_seg_0:reset_n, seven_seg_1:reset_n, seven_seg_2:reset_n, seven_seg_3:reset_n, seven_seg_4:reset_n, seven_seg_5:reset_n, switches:reset_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [NIOSII:reset_req, SDRAM:reset_req, rst_translator:reset_req_in]
	wire         niosii_debug_reset_request_reset;                                 // NIOSII:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [JTAG:rst_n, mm_interconnect_0:JTAG_reset_reset_bridge_in_reset_reset]

	System_Audio_Video audio_video (
		.clk         (clk_clk),                                                          //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                   //                  reset.reset
		.address     (mm_interconnect_0_audio_video_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_video_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_video_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_video_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_video_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_video_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_video_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (aud_vid_SDAT),                                                     //     external_interface.export
		.I2C_SCLK    (aud_vid_SCLK)                                                      //                       .export
	);

	System_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	System_NIOSII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (niosii_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosii_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	System_SDRAM sdram (
		.clk        (clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_sdram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sdram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sdram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sdram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sdram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sdram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sdram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	System_Timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	System_key_0 key_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_0_s1_readdata),   //                    .readdata
		.in_port    (key_0_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)               //                 irq.irq
	);

	System_key_0 key_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_1_s1_readdata),   //                    .readdata
		.in_port    (key_1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)               //                 irq.irq
	);

	System_key_0 key_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_2_s1_readdata),   //                    .readdata
		.in_port    (key_2_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)               //                 irq.irq
	);

	System_key_0 key_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_3_s1_readdata),   //                    .readdata
		.in_port    (key_3_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)               //                 irq.irq
	);

	System_red_leds red_leds (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_red_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_leds_s1_readdata),   //                    .readdata
		.out_port   (red_leds_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_0_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_0_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_2_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_2_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_3_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_3_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_4_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_4_export)                           // external_connection.export
	);

	System_seven_seg_0 seven_seg_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_5_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_5_export)                           // external_connection.export
	);

	System_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	System_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                          //                          clk_0_clk.clk
		.JTAG_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                               //   JTAG_reset_reset_bridge_in_reset.reset
		.NIOSII_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                   // NIOSII_reset_reset_bridge_in_reset.reset
		.NIOSII_data_master_address                     (niosii_data_master_address),                                       //                 NIOSII_data_master.address
		.NIOSII_data_master_waitrequest                 (niosii_data_master_waitrequest),                                   //                                   .waitrequest
		.NIOSII_data_master_byteenable                  (niosii_data_master_byteenable),                                    //                                   .byteenable
		.NIOSII_data_master_read                        (niosii_data_master_read),                                          //                                   .read
		.NIOSII_data_master_readdata                    (niosii_data_master_readdata),                                      //                                   .readdata
		.NIOSII_data_master_readdatavalid               (niosii_data_master_readdatavalid),                                 //                                   .readdatavalid
		.NIOSII_data_master_write                       (niosii_data_master_write),                                         //                                   .write
		.NIOSII_data_master_writedata                   (niosii_data_master_writedata),                                     //                                   .writedata
		.NIOSII_data_master_debugaccess                 (niosii_data_master_debugaccess),                                   //                                   .debugaccess
		.NIOSII_instruction_master_address              (niosii_instruction_master_address),                                //          NIOSII_instruction_master.address
		.NIOSII_instruction_master_waitrequest          (niosii_instruction_master_waitrequest),                            //                                   .waitrequest
		.NIOSII_instruction_master_read                 (niosii_instruction_master_read),                                   //                                   .read
		.NIOSII_instruction_master_readdata             (niosii_instruction_master_readdata),                               //                                   .readdata
		.NIOSII_instruction_master_readdatavalid        (niosii_instruction_master_readdatavalid),                          //                                   .readdatavalid
		.Audio_Video_avalon_av_config_slave_address     (mm_interconnect_0_audio_video_avalon_av_config_slave_address),     // Audio_Video_avalon_av_config_slave.address
		.Audio_Video_avalon_av_config_slave_write       (mm_interconnect_0_audio_video_avalon_av_config_slave_write),       //                                   .write
		.Audio_Video_avalon_av_config_slave_read        (mm_interconnect_0_audio_video_avalon_av_config_slave_read),        //                                   .read
		.Audio_Video_avalon_av_config_slave_readdata    (mm_interconnect_0_audio_video_avalon_av_config_slave_readdata),    //                                   .readdata
		.Audio_Video_avalon_av_config_slave_writedata   (mm_interconnect_0_audio_video_avalon_av_config_slave_writedata),   //                                   .writedata
		.Audio_Video_avalon_av_config_slave_byteenable  (mm_interconnect_0_audio_video_avalon_av_config_slave_byteenable),  //                                   .byteenable
		.Audio_Video_avalon_av_config_slave_waitrequest (mm_interconnect_0_audio_video_avalon_av_config_slave_waitrequest), //                                   .waitrequest
		.JTAG_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_avalon_jtag_slave_address),                 //             JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_avalon_jtag_slave_write),                   //                                   .write
		.JTAG_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_avalon_jtag_slave_read),                    //                                   .read
		.JTAG_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                //                                   .readdata
		.JTAG_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),               //                                   .writedata
		.JTAG_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),             //                                   .waitrequest
		.JTAG_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),              //                                   .chipselect
		.key_0_s1_address                               (mm_interconnect_0_key_0_s1_address),                               //                           key_0_s1.address
		.key_0_s1_write                                 (mm_interconnect_0_key_0_s1_write),                                 //                                   .write
		.key_0_s1_readdata                              (mm_interconnect_0_key_0_s1_readdata),                              //                                   .readdata
		.key_0_s1_writedata                             (mm_interconnect_0_key_0_s1_writedata),                             //                                   .writedata
		.key_0_s1_chipselect                            (mm_interconnect_0_key_0_s1_chipselect),                            //                                   .chipselect
		.key_1_s1_address                               (mm_interconnect_0_key_1_s1_address),                               //                           key_1_s1.address
		.key_1_s1_write                                 (mm_interconnect_0_key_1_s1_write),                                 //                                   .write
		.key_1_s1_readdata                              (mm_interconnect_0_key_1_s1_readdata),                              //                                   .readdata
		.key_1_s1_writedata                             (mm_interconnect_0_key_1_s1_writedata),                             //                                   .writedata
		.key_1_s1_chipselect                            (mm_interconnect_0_key_1_s1_chipselect),                            //                                   .chipselect
		.key_2_s1_address                               (mm_interconnect_0_key_2_s1_address),                               //                           key_2_s1.address
		.key_2_s1_write                                 (mm_interconnect_0_key_2_s1_write),                                 //                                   .write
		.key_2_s1_readdata                              (mm_interconnect_0_key_2_s1_readdata),                              //                                   .readdata
		.key_2_s1_writedata                             (mm_interconnect_0_key_2_s1_writedata),                             //                                   .writedata
		.key_2_s1_chipselect                            (mm_interconnect_0_key_2_s1_chipselect),                            //                                   .chipselect
		.key_3_s1_address                               (mm_interconnect_0_key_3_s1_address),                               //                           key_3_s1.address
		.key_3_s1_write                                 (mm_interconnect_0_key_3_s1_write),                                 //                                   .write
		.key_3_s1_readdata                              (mm_interconnect_0_key_3_s1_readdata),                              //                                   .readdata
		.key_3_s1_writedata                             (mm_interconnect_0_key_3_s1_writedata),                             //                                   .writedata
		.key_3_s1_chipselect                            (mm_interconnect_0_key_3_s1_chipselect),                            //                                   .chipselect
		.NIOSII_debug_mem_slave_address                 (mm_interconnect_0_niosii_debug_mem_slave_address),                 //             NIOSII_debug_mem_slave.address
		.NIOSII_debug_mem_slave_write                   (mm_interconnect_0_niosii_debug_mem_slave_write),                   //                                   .write
		.NIOSII_debug_mem_slave_read                    (mm_interconnect_0_niosii_debug_mem_slave_read),                    //                                   .read
		.NIOSII_debug_mem_slave_readdata                (mm_interconnect_0_niosii_debug_mem_slave_readdata),                //                                   .readdata
		.NIOSII_debug_mem_slave_writedata               (mm_interconnect_0_niosii_debug_mem_slave_writedata),               //                                   .writedata
		.NIOSII_debug_mem_slave_byteenable              (mm_interconnect_0_niosii_debug_mem_slave_byteenable),              //                                   .byteenable
		.NIOSII_debug_mem_slave_waitrequest             (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),             //                                   .waitrequest
		.NIOSII_debug_mem_slave_debugaccess             (mm_interconnect_0_niosii_debug_mem_slave_debugaccess),             //                                   .debugaccess
		.red_leds_s1_address                            (mm_interconnect_0_red_leds_s1_address),                            //                        red_leds_s1.address
		.red_leds_s1_write                              (mm_interconnect_0_red_leds_s1_write),                              //                                   .write
		.red_leds_s1_readdata                           (mm_interconnect_0_red_leds_s1_readdata),                           //                                   .readdata
		.red_leds_s1_writedata                          (mm_interconnect_0_red_leds_s1_writedata),                          //                                   .writedata
		.red_leds_s1_chipselect                         (mm_interconnect_0_red_leds_s1_chipselect),                         //                                   .chipselect
		.SDRAM_s1_address                               (mm_interconnect_0_sdram_s1_address),                               //                           SDRAM_s1.address
		.SDRAM_s1_write                                 (mm_interconnect_0_sdram_s1_write),                                 //                                   .write
		.SDRAM_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                              //                                   .readdata
		.SDRAM_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                             //                                   .writedata
		.SDRAM_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                            //                                   .byteenable
		.SDRAM_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                            //                                   .chipselect
		.SDRAM_s1_clken                                 (mm_interconnect_0_sdram_s1_clken),                                 //                                   .clken
		.seven_seg_0_s1_address                         (mm_interconnect_0_seven_seg_0_s1_address),                         //                     seven_seg_0_s1.address
		.seven_seg_0_s1_write                           (mm_interconnect_0_seven_seg_0_s1_write),                           //                                   .write
		.seven_seg_0_s1_readdata                        (mm_interconnect_0_seven_seg_0_s1_readdata),                        //                                   .readdata
		.seven_seg_0_s1_writedata                       (mm_interconnect_0_seven_seg_0_s1_writedata),                       //                                   .writedata
		.seven_seg_0_s1_chipselect                      (mm_interconnect_0_seven_seg_0_s1_chipselect),                      //                                   .chipselect
		.seven_seg_1_s1_address                         (mm_interconnect_0_seven_seg_1_s1_address),                         //                     seven_seg_1_s1.address
		.seven_seg_1_s1_write                           (mm_interconnect_0_seven_seg_1_s1_write),                           //                                   .write
		.seven_seg_1_s1_readdata                        (mm_interconnect_0_seven_seg_1_s1_readdata),                        //                                   .readdata
		.seven_seg_1_s1_writedata                       (mm_interconnect_0_seven_seg_1_s1_writedata),                       //                                   .writedata
		.seven_seg_1_s1_chipselect                      (mm_interconnect_0_seven_seg_1_s1_chipselect),                      //                                   .chipselect
		.seven_seg_2_s1_address                         (mm_interconnect_0_seven_seg_2_s1_address),                         //                     seven_seg_2_s1.address
		.seven_seg_2_s1_write                           (mm_interconnect_0_seven_seg_2_s1_write),                           //                                   .write
		.seven_seg_2_s1_readdata                        (mm_interconnect_0_seven_seg_2_s1_readdata),                        //                                   .readdata
		.seven_seg_2_s1_writedata                       (mm_interconnect_0_seven_seg_2_s1_writedata),                       //                                   .writedata
		.seven_seg_2_s1_chipselect                      (mm_interconnect_0_seven_seg_2_s1_chipselect),                      //                                   .chipselect
		.seven_seg_3_s1_address                         (mm_interconnect_0_seven_seg_3_s1_address),                         //                     seven_seg_3_s1.address
		.seven_seg_3_s1_write                           (mm_interconnect_0_seven_seg_3_s1_write),                           //                                   .write
		.seven_seg_3_s1_readdata                        (mm_interconnect_0_seven_seg_3_s1_readdata),                        //                                   .readdata
		.seven_seg_3_s1_writedata                       (mm_interconnect_0_seven_seg_3_s1_writedata),                       //                                   .writedata
		.seven_seg_3_s1_chipselect                      (mm_interconnect_0_seven_seg_3_s1_chipselect),                      //                                   .chipselect
		.seven_seg_4_s1_address                         (mm_interconnect_0_seven_seg_4_s1_address),                         //                     seven_seg_4_s1.address
		.seven_seg_4_s1_write                           (mm_interconnect_0_seven_seg_4_s1_write),                           //                                   .write
		.seven_seg_4_s1_readdata                        (mm_interconnect_0_seven_seg_4_s1_readdata),                        //                                   .readdata
		.seven_seg_4_s1_writedata                       (mm_interconnect_0_seven_seg_4_s1_writedata),                       //                                   .writedata
		.seven_seg_4_s1_chipselect                      (mm_interconnect_0_seven_seg_4_s1_chipselect),                      //                                   .chipselect
		.seven_seg_5_s1_address                         (mm_interconnect_0_seven_seg_5_s1_address),                         //                     seven_seg_5_s1.address
		.seven_seg_5_s1_write                           (mm_interconnect_0_seven_seg_5_s1_write),                           //                                   .write
		.seven_seg_5_s1_readdata                        (mm_interconnect_0_seven_seg_5_s1_readdata),                        //                                   .readdata
		.seven_seg_5_s1_writedata                       (mm_interconnect_0_seven_seg_5_s1_writedata),                       //                                   .writedata
		.seven_seg_5_s1_chipselect                      (mm_interconnect_0_seven_seg_5_s1_chipselect),                      //                                   .chipselect
		.switches_s1_address                            (mm_interconnect_0_switches_s1_address),                            //                        switches_s1.address
		.switches_s1_readdata                           (mm_interconnect_0_switches_s1_readdata),                           //                                   .readdata
		.Timer_s1_address                               (mm_interconnect_0_timer_s1_address),                               //                           Timer_s1.address
		.Timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                                 //                                   .write
		.Timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                              //                                   .readdata
		.Timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                             //                                   .writedata
		.Timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect)                             //                                   .chipselect
	);

	System_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (niosii_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (niosii_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
