// test.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module test (
		input  wire        audio_ADCDAT,    //     audio.ADCDAT
		input  wire        audio_ADCLRCK,   //          .ADCLRCK
		input  wire        audio_BCLK,      //          .BCLK
		output wire        audio_DACDAT,    //          .DACDAT
		input  wire        audio_DACLRCK,   //          .DACLRCK
		output wire        audio_clk_clk,   // audio_clk.clk
		input  wire        button_1_export, //  button_1.export
		input  wire        button_2_export, //  button_2.export
		input  wire        clk_clk,         //       clk.clk
		input  wire        reset_reset_n,   //     reset.reset_n
		input  wire        rs232_RXD,       //     rs232.RXD
		output wire        rs232_TXD,       //          .TXD
		output wire [12:0] sdram_addr,      //     sdram.addr
		output wire [1:0]  sdram_ba,        //          .ba
		output wire        sdram_cas_n,     //          .cas_n
		output wire        sdram_cke,       //          .cke
		output wire        sdram_cs_n,      //          .cs_n
		inout  wire [15:0] sdram_dq,        //          .dq
		output wire [1:0]  sdram_dqm,       //          .dqm
		output wire        sdram_ras_n,     //          .ras_n
		output wire        sdram_we_n,      //          .we_n
		output wire        sdram_clk_clk,   // sdram_clk.clk
		output wire        vga_CLK,         //       vga.CLK
		output wire        vga_HS,          //          .HS
		output wire        vga_VS,          //          .VS
		output wire        vga_BLANK,       //          .BLANK
		output wire        vga_SYNC,        //          .SYNC
		output wire [7:0]  vga_R,           //          .R
		output wire [7:0]  vga_G,           //          .G
		output wire [7:0]  vga_B            //          .B
	);

	wire         alpha_blender_avalon_blended_source_valid;                          // Alpha_Blender:output_valid -> Dual_Clock_FIFO:stream_in_valid
	wire  [29:0] alpha_blender_avalon_blended_source_data;                           // Alpha_Blender:output_data -> Dual_Clock_FIFO:stream_in_data
	wire         alpha_blender_avalon_blended_source_ready;                          // Dual_Clock_FIFO:stream_in_ready -> Alpha_Blender:output_ready
	wire         alpha_blender_avalon_blended_source_startofpacket;                  // Alpha_Blender:output_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	wire         alpha_blender_avalon_blended_source_endofpacket;                    // Alpha_Blender:output_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	wire         char_buffer_avalon_char_source_valid;                               // Char_Buffer:stream_valid -> Alpha_Blender:foreground_valid
	wire  [39:0] char_buffer_avalon_char_source_data;                                // Char_Buffer:stream_data -> Alpha_Blender:foreground_data
	wire         char_buffer_avalon_char_source_ready;                               // Alpha_Blender:foreground_ready -> Char_Buffer:stream_ready
	wire         char_buffer_avalon_char_source_startofpacket;                       // Char_Buffer:stream_startofpacket -> Alpha_Blender:foreground_startofpacket
	wire         char_buffer_avalon_char_source_endofpacket;                         // Char_Buffer:stream_endofpacket -> Alpha_Blender:foreground_endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                      // Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                       // Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                      // VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;              // Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                // Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         pixel_buffer_avalon_pixel_source_valid;                             // Pixel_Buffer:stream_valid -> RGB_Resampler:stream_in_valid
	wire   [7:0] pixel_buffer_avalon_pixel_source_data;                              // Pixel_Buffer:stream_data -> RGB_Resampler:stream_in_data
	wire         pixel_buffer_avalon_pixel_source_ready;                             // RGB_Resampler:stream_in_ready -> Pixel_Buffer:stream_ready
	wire         pixel_buffer_avalon_pixel_source_startofpacket;                     // Pixel_Buffer:stream_startofpacket -> RGB_Resampler:stream_in_startofpacket
	wire         pixel_buffer_avalon_pixel_source_endofpacket;                       // Pixel_Buffer:stream_endofpacket -> RGB_Resampler:stream_in_endofpacket
	wire         rgb_resampler_avalon_rgb_source_valid;                              // RGB_Resampler:stream_out_valid -> Alpha_Blender:background_valid
	wire  [29:0] rgb_resampler_avalon_rgb_source_data;                               // RGB_Resampler:stream_out_data -> Alpha_Blender:background_data
	wire         rgb_resampler_avalon_rgb_source_ready;                              // Alpha_Blender:background_ready -> RGB_Resampler:stream_out_ready
	wire         rgb_resampler_avalon_rgb_source_startofpacket;                      // RGB_Resampler:stream_out_startofpacket -> Alpha_Blender:background_startofpacket
	wire         rgb_resampler_avalon_rgb_source_endofpacket;                        // RGB_Resampler:stream_out_endofpacket -> Alpha_Blender:background_endofpacket
	wire         sys_clk_sys_clk_clk;                                                // Sys_Clk:sys_clk_clk -> [Alpha_Blender:clk, Audio:clk, Audio_Clk:ref_clk_clk, CPU:clk, Char_Buffer:clk, Dual_Clock_FIFO:clk_stream_in, JTAG:clk, Onchip_Memory:clk, Pixel_Buffer:clk, RGB_Resampler:clk, SDRAM:clk, Video_Clk:ref_clk_clk, WIFI_Serial_Port:clk, button_1:clk, button_2:clk, irq_mapper:clk, mm_interconnect_0:Sys_Clk_sys_clk_clk, rst_controller:clk, rst_controller_002:clk, timer:clk, timer_0:clk]
	wire         video_clk_vga_clk_clk;                                              // Video_Clk:vga_clk_clk -> [Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_001:clk, rst_controller_004:clk]
	wire         sys_clk_reset_source_reset;                                         // Sys_Clk:reset_source_reset -> [Audio_Clk:ref_reset_reset, rst_controller_005:reset_in1]
	wire         pixel_buffer_avalon_pixel_dma_master_waitrequest;                   // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_waitrequest -> Pixel_Buffer:master_waitrequest
	wire   [7:0] pixel_buffer_avalon_pixel_dma_master_readdata;                      // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_readdata -> Pixel_Buffer:master_readdata
	wire  [31:0] pixel_buffer_avalon_pixel_dma_master_address;                       // Pixel_Buffer:master_address -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_address
	wire         pixel_buffer_avalon_pixel_dma_master_read;                          // Pixel_Buffer:master_read -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_read
	wire         pixel_buffer_avalon_pixel_dma_master_readdatavalid;                 // mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_readdatavalid -> Pixel_Buffer:master_readdatavalid
	wire         pixel_buffer_avalon_pixel_dma_master_lock;                          // Pixel_Buffer:master_arbiterlock -> mm_interconnect_0:Pixel_Buffer_avalon_pixel_dma_master_lock
	wire  [31:0] cpu_data_master_readdata;                                           // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                                        // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                                        // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                            // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                         // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                               // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_readdatavalid;                                      // mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	wire         cpu_data_master_write;                                              // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                          // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                    // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                                 // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                     // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                        // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                               // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;              // mm_interconnect_0:Audio_avalon_audio_slave_chipselect -> Audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;                // Audio:readdata -> mm_interconnect_0:Audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                 // mm_interconnect_0:Audio_avalon_audio_slave_address -> Audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                    // mm_interconnect_0:Audio_avalon_audio_slave_read -> Audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                   // mm_interconnect_0:Audio_avalon_audio_slave_write -> Audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;               // mm_interconnect_0:Audio_avalon_audio_slave_writedata -> Audio:writedata
	wire         mm_interconnect_0_char_buffer_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_chipselect -> Char_Buffer:buf_chipselect
	wire   [7:0] mm_interconnect_0_char_buffer_avalon_char_buffer_slave_readdata;    // Char_Buffer:buf_readdata -> mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_char_buffer_avalon_char_buffer_slave_waitrequest; // Char_Buffer:buf_waitrequest -> mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_char_buffer_avalon_char_buffer_slave_address;     // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_address -> Char_Buffer:buf_address
	wire         mm_interconnect_0_char_buffer_avalon_char_buffer_slave_read;        // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_read -> Char_Buffer:buf_read
	wire   [0:0] mm_interconnect_0_char_buffer_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_byteenable -> Char_Buffer:buf_byteenable
	wire         mm_interconnect_0_char_buffer_avalon_char_buffer_slave_write;       // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_write -> Char_Buffer:buf_write
	wire   [7:0] mm_interconnect_0_char_buffer_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:Char_Buffer_avalon_char_buffer_slave_writedata -> Char_Buffer:buf_writedata
	wire         mm_interconnect_0_char_buffer_avalon_char_control_slave_chipselect; // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_chipselect -> Char_Buffer:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_char_buffer_avalon_char_control_slave_readdata;   // Char_Buffer:ctrl_readdata -> mm_interconnect_0:Char_Buffer_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_char_buffer_avalon_char_control_slave_address;    // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_address -> Char_Buffer:ctrl_address
	wire         mm_interconnect_0_char_buffer_avalon_char_control_slave_read;       // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_read -> Char_Buffer:ctrl_read
	wire   [3:0] mm_interconnect_0_char_buffer_avalon_char_control_slave_byteenable; // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_byteenable -> Char_Buffer:ctrl_byteenable
	wire         mm_interconnect_0_char_buffer_avalon_char_control_slave_write;      // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_write -> Char_Buffer:ctrl_write
	wire  [31:0] mm_interconnect_0_char_buffer_avalon_char_control_slave_writedata;  // mm_interconnect_0:Char_Buffer_avalon_char_control_slave_writedata -> Char_Buffer:ctrl_writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata;       // Pixel_Buffer:slave_readdata -> mm_interconnect_0:Pixel_Buffer_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_address;        // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_address -> Pixel_Buffer:slave_address
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_read;           // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_read -> Pixel_Buffer:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable;     // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_byteenable -> Pixel_Buffer:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_avalon_control_slave_write;          // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_write -> Pixel_Buffer:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata;      // mm_interconnect_0:Pixel_Buffer_avalon_control_slave_writedata -> Pixel_Buffer:slave_writedata
	wire  [31:0] mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata;          // RGB_Resampler:slave_readdata -> mm_interconnect_0:RGB_Resampler_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read;              // mm_interconnect_0:RGB_Resampler_avalon_rgb_slave_read -> RGB_Resampler:slave_read
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                     // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                  // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                  // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                      // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                         // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                   // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                        // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                    // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                      // mm_interconnect_0:Onchip_Memory_s1_chipselect -> Onchip_Memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                        // Onchip_Memory:readdata -> mm_interconnect_0:Onchip_Memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                         // mm_interconnect_0:Onchip_Memory_s1_address -> Onchip_Memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                      // mm_interconnect_0:Onchip_Memory_s1_byteenable -> Onchip_Memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                           // mm_interconnect_0:Onchip_Memory_s1_write -> Onchip_Memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                       // mm_interconnect_0:Onchip_Memory_s1_writedata -> Onchip_Memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                           // mm_interconnect_0:Onchip_Memory_s1_clken -> Onchip_Memory:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                  // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;               // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                   // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                      // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                     // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                 // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire         mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_chipselect;   // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_chipselect -> WIFI_Serial_Port:chipselect
	wire  [31:0] mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_readdata;     // WIFI_Serial_Port:readdata -> mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_address;      // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_address -> WIFI_Serial_Port:address
	wire         mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_read;         // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_read -> WIFI_Serial_Port:read
	wire   [3:0] mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_byteenable;   // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_byteenable -> WIFI_Serial_Port:byteenable
	wire         mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_write;        // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_write -> WIFI_Serial_Port:write
	wire  [31:0] mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_writedata;    // mm_interconnect_0:WIFI_Serial_Port_avalon_rs232_slave_writedata -> WIFI_Serial_Port:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                            // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                              // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                               // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                 // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                             // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_button_1_s1_chipselect;                           // mm_interconnect_0:button_1_s1_chipselect -> button_1:chipselect
	wire  [31:0] mm_interconnect_0_button_1_s1_readdata;                             // button_1:readdata -> mm_interconnect_0:button_1_s1_readdata
	wire   [1:0] mm_interconnect_0_button_1_s1_address;                              // mm_interconnect_0:button_1_s1_address -> button_1:address
	wire         mm_interconnect_0_button_1_s1_write;                                // mm_interconnect_0:button_1_s1_write -> button_1:write_n
	wire  [31:0] mm_interconnect_0_button_1_s1_writedata;                            // mm_interconnect_0:button_1_s1_writedata -> button_1:writedata
	wire         mm_interconnect_0_button_2_s1_chipselect;                           // mm_interconnect_0:button_2_s1_chipselect -> button_2:chipselect
	wire  [31:0] mm_interconnect_0_button_2_s1_readdata;                             // button_2:readdata -> mm_interconnect_0:button_2_s1_readdata
	wire   [1:0] mm_interconnect_0_button_2_s1_address;                              // mm_interconnect_0:button_2_s1_address -> button_2:address
	wire         mm_interconnect_0_button_2_s1_write;                                // mm_interconnect_0:button_2_s1_write -> button_2:write_n
	wire  [31:0] mm_interconnect_0_button_2_s1_writedata;                            // mm_interconnect_0:button_2_s1_writedata -> button_2:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                              // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                 // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                   // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                               // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         irq_mapper_receiver0_irq;                                           // Audio:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // WIFI_Serial_Port:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // JTAG:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                           // button_2:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                           // button_1:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                           // timer:irq -> irq_mapper:receiver6_irq
	wire  [31:0] cpu_irq_irq;                                                        // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Alpha_Blender:reset, Audio:reset, CPU:reset_n, Char_Buffer:reset, Dual_Clock_FIFO:reset_stream_in, Onchip_Memory:reset, Pixel_Buffer:reset, RGB_Resampler:reset, SDRAM:reset_n, irq_mapper:reset, mm_interconnect_0:Pixel_Buffer_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [CPU:reset_req, Onchip_Memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                      // CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in0]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> Dual_Clock_FIFO:reset_stream_out
	wire         rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [JTAG:rst_n, WIFI_Serial_Port:reset, button_1:reset_n, button_2:reset_n, mm_interconnect_0:JTAG_reset_reset_bridge_in_reset_reset, timer:reset_n, timer_0:reset_n]
	wire         rst_controller_003_reset_out_reset;                                 // rst_controller_003:reset_out -> Sys_Clk:ref_reset_reset
	wire         rst_controller_004_reset_out_reset;                                 // rst_controller_004:reset_out -> VGA_Controller:reset
	wire         video_clk_reset_source_reset;                                       // Video_Clk:reset_source_reset -> rst_controller_004:reset_in2
	wire         rst_controller_005_reset_out_reset;                                 // rst_controller_005:reset_out -> Video_Clk:ref_reset_reset

	test_Alpha_Blender alpha_blender (
		.clk                      (sys_clk_sys_clk_clk),                               //                    clk.clk
		.reset                    (rst_controller_reset_out_reset),                    //                  reset.reset
		.foreground_data          (char_buffer_avalon_char_source_data),               // avalon_foreground_sink.data
		.foreground_startofpacket (char_buffer_avalon_char_source_startofpacket),      //                       .startofpacket
		.foreground_endofpacket   (char_buffer_avalon_char_source_endofpacket),        //                       .endofpacket
		.foreground_valid         (char_buffer_avalon_char_source_valid),              //                       .valid
		.foreground_ready         (char_buffer_avalon_char_source_ready),              //                       .ready
		.background_data          (rgb_resampler_avalon_rgb_source_data),              // avalon_background_sink.data
		.background_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),     //                       .startofpacket
		.background_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),       //                       .endofpacket
		.background_valid         (rgb_resampler_avalon_rgb_source_valid),             //                       .valid
		.background_ready         (rgb_resampler_avalon_rgb_source_ready),             //                       .ready
		.output_ready             (alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	test_Audio audio (
		.clk         (sys_clk_sys_clk_clk),                                   //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                              //          interrupt.irq
		.AUD_ADCDAT  (audio_ADCDAT),                                          // external_interface.export
		.AUD_ADCLRCK (audio_ADCLRCK),                                         //                   .export
		.AUD_BCLK    (audio_BCLK),                                            //                   .export
		.AUD_DACDAT  (audio_DACDAT),                                          //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                          //                   .export
	);

	test_Audio_Clk audio_clk (
		.ref_clk_clk        (sys_clk_sys_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (sys_clk_reset_source_reset), //    ref_reset.reset
		.audio_clk_clk      (audio_clk_clk),              //    audio_clk.clk
		.reset_source_reset ()                            // reset_source.reset
	);

	test_CPU cpu (
		.clk                                 (sys_clk_sys_clk_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	test_Char_Buffer char_buffer (
		.clk                  (sys_clk_sys_clk_clk),                                                //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                     //                     reset.reset
		.ctrl_address         (mm_interconnect_0_char_buffer_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_char_buffer_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_char_buffer_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_char_buffer_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_char_buffer_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_char_buffer_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_char_buffer_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (char_buffer_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (char_buffer_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (char_buffer_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (char_buffer_avalon_char_source_valid),                               //                          .valid
		.stream_data          (char_buffer_avalon_char_source_data)                                 //                          .data
	);

	test_Dual_Clock_FIFO dual_clock_fifo (
		.clk_stream_in            (sys_clk_sys_clk_clk),                                   //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                        //         reset_stream_in.reset
		.clk_stream_out           (video_clk_vga_clk_clk),                                 //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                    //        reset_stream_out.reset
		.stream_in_ready          (alpha_blender_avalon_blended_source_ready),             //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blender_avalon_blended_source_startofpacket),     //                        .startofpacket
		.stream_in_endofpacket    (alpha_blender_avalon_blended_source_endofpacket),       //                        .endofpacket
		.stream_in_valid          (alpha_blender_avalon_blended_source_valid),             //                        .valid
		.stream_in_data           (alpha_blender_avalon_blended_source_data),              //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	test_JTAG jtag (
		.clk            (sys_clk_sys_clk_clk),                                  //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                              //               irq.irq
	);

	test_Onchip_Memory onchip_memory (
		.clk        (sys_clk_sys_clk_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	test_Pixel_Buffer pixel_buffer (
		.clk                  (sys_clk_sys_clk_clk),                                            //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                 //                   reset.reset
		.master_readdatavalid (pixel_buffer_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_avalon_pixel_source_data)                           //                        .data
	);

	test_RGB_Resampler rgb_resampler (
		.clk                      (sys_clk_sys_clk_clk),                                       //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                            //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_avalon_pixel_source_startofpacket),            //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_avalon_pixel_source_endofpacket),              //                  .endofpacket
		.stream_in_valid          (pixel_buffer_avalon_pixel_source_valid),                    //                  .valid
		.stream_in_ready          (pixel_buffer_avalon_pixel_source_ready),                    //                  .ready
		.stream_in_data           (pixel_buffer_avalon_pixel_source_data),                     //                  .data
		.slave_read               (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                       //                  .data
	);

	test_SDRAM sdram (
		.clk            (sys_clk_sys_clk_clk),                      //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	test_Sys_Clk sys_clk (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_clk_sys_clk_clk),                //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_clk_reset_source_reset)          // reset_source.reset
	);

	test_VGA_Controller vga_controller (
		.clk           (video_clk_vga_clk_clk),                                 //                clk.clk
		.reset         (rst_controller_004_reset_out_reset),                    //              reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                               // external_interface.export
		.VGA_HS        (vga_HS),                                                //                   .export
		.VGA_VS        (vga_VS),                                                //                   .export
		.VGA_BLANK     (vga_BLANK),                                             //                   .export
		.VGA_SYNC      (vga_SYNC),                                              //                   .export
		.VGA_R         (vga_R),                                                 //                   .export
		.VGA_G         (vga_G),                                                 //                   .export
		.VGA_B         (vga_B)                                                  //                   .export
	);

	test_Video_Clk video_clk (
		.ref_clk_clk        (sys_clk_sys_clk_clk),                //      ref_clk.clk
		.ref_reset_reset    (rst_controller_005_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_clk_vga_clk_clk),              //      vga_clk.clk
		.reset_source_reset (video_clk_reset_source_reset)        // reset_source.reset
	);

	test_WIFI_Serial_Port wifi_serial_port (
		.clk        (sys_clk_sys_clk_clk),                                              //                clk.clk
		.reset      (rst_controller_002_reset_out_reset),                               //              reset.reset
		.address    (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver1_irq),                                         //          interrupt.irq
		.UART_RXD   (rs232_RXD),                                                        // external_interface.export
		.UART_TXD   (rs232_TXD)                                                         //                   .export
	);

	test_button_1 button_1 (
		.clk        (sys_clk_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_button_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_1_s1_readdata),   //                    .readdata
		.in_port    (button_1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                  //                 irq.irq
	);

	test_button_1 button_2 (
		.clk        (sys_clk_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_button_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_2_s1_readdata),   //                    .readdata
		.in_port    (button_2_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                  //                 irq.irq
	);

	test_timer timer (
		.clk        (sys_clk_sys_clk_clk),                   //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)               //   irq.irq
	);

	test_timer timer_0 (
		.clk        (sys_clk_sys_clk_clk),                     //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	test_mm_interconnect_0 mm_interconnect_0 (
		.Sys_Clk_sys_clk_clk                                (sys_clk_sys_clk_clk),                                                //                          Sys_Clk_sys_clk.clk
		.JTAG_reset_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                                 //         JTAG_reset_reset_bridge_in_reset.reset
		.Pixel_Buffer_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                     // Pixel_Buffer_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                            (cpu_data_master_address),                                            //                          CPU_data_master.address
		.CPU_data_master_waitrequest                        (cpu_data_master_waitrequest),                                        //                                         .waitrequest
		.CPU_data_master_byteenable                         (cpu_data_master_byteenable),                                         //                                         .byteenable
		.CPU_data_master_read                               (cpu_data_master_read),                                               //                                         .read
		.CPU_data_master_readdata                           (cpu_data_master_readdata),                                           //                                         .readdata
		.CPU_data_master_readdatavalid                      (cpu_data_master_readdatavalid),                                      //                                         .readdatavalid
		.CPU_data_master_write                              (cpu_data_master_write),                                              //                                         .write
		.CPU_data_master_writedata                          (cpu_data_master_writedata),                                          //                                         .writedata
		.CPU_data_master_debugaccess                        (cpu_data_master_debugaccess),                                        //                                         .debugaccess
		.CPU_instruction_master_address                     (cpu_instruction_master_address),                                     //                   CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                 (cpu_instruction_master_waitrequest),                                 //                                         .waitrequest
		.CPU_instruction_master_read                        (cpu_instruction_master_read),                                        //                                         .read
		.CPU_instruction_master_readdata                    (cpu_instruction_master_readdata),                                    //                                         .readdata
		.CPU_instruction_master_readdatavalid               (cpu_instruction_master_readdatavalid),                               //                                         .readdatavalid
		.Pixel_Buffer_avalon_pixel_dma_master_address       (pixel_buffer_avalon_pixel_dma_master_address),                       //     Pixel_Buffer_avalon_pixel_dma_master.address
		.Pixel_Buffer_avalon_pixel_dma_master_waitrequest   (pixel_buffer_avalon_pixel_dma_master_waitrequest),                   //                                         .waitrequest
		.Pixel_Buffer_avalon_pixel_dma_master_read          (pixel_buffer_avalon_pixel_dma_master_read),                          //                                         .read
		.Pixel_Buffer_avalon_pixel_dma_master_readdata      (pixel_buffer_avalon_pixel_dma_master_readdata),                      //                                         .readdata
		.Pixel_Buffer_avalon_pixel_dma_master_readdatavalid (pixel_buffer_avalon_pixel_dma_master_readdatavalid),                 //                                         .readdatavalid
		.Pixel_Buffer_avalon_pixel_dma_master_lock          (pixel_buffer_avalon_pixel_dma_master_lock),                          //                                         .lock
		.Audio_avalon_audio_slave_address                   (mm_interconnect_0_audio_avalon_audio_slave_address),                 //                 Audio_avalon_audio_slave.address
		.Audio_avalon_audio_slave_write                     (mm_interconnect_0_audio_avalon_audio_slave_write),                   //                                         .write
		.Audio_avalon_audio_slave_read                      (mm_interconnect_0_audio_avalon_audio_slave_read),                    //                                         .read
		.Audio_avalon_audio_slave_readdata                  (mm_interconnect_0_audio_avalon_audio_slave_readdata),                //                                         .readdata
		.Audio_avalon_audio_slave_writedata                 (mm_interconnect_0_audio_avalon_audio_slave_writedata),               //                                         .writedata
		.Audio_avalon_audio_slave_chipselect                (mm_interconnect_0_audio_avalon_audio_slave_chipselect),              //                                         .chipselect
		.button_1_s1_address                                (mm_interconnect_0_button_1_s1_address),                              //                              button_1_s1.address
		.button_1_s1_write                                  (mm_interconnect_0_button_1_s1_write),                                //                                         .write
		.button_1_s1_readdata                               (mm_interconnect_0_button_1_s1_readdata),                             //                                         .readdata
		.button_1_s1_writedata                              (mm_interconnect_0_button_1_s1_writedata),                            //                                         .writedata
		.button_1_s1_chipselect                             (mm_interconnect_0_button_1_s1_chipselect),                           //                                         .chipselect
		.button_2_s1_address                                (mm_interconnect_0_button_2_s1_address),                              //                              button_2_s1.address
		.button_2_s1_write                                  (mm_interconnect_0_button_2_s1_write),                                //                                         .write
		.button_2_s1_readdata                               (mm_interconnect_0_button_2_s1_readdata),                             //                                         .readdata
		.button_2_s1_writedata                              (mm_interconnect_0_button_2_s1_writedata),                            //                                         .writedata
		.button_2_s1_chipselect                             (mm_interconnect_0_button_2_s1_chipselect),                           //                                         .chipselect
		.Char_Buffer_avalon_char_buffer_slave_address       (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_address),     //     Char_Buffer_avalon_char_buffer_slave.address
		.Char_Buffer_avalon_char_buffer_slave_write         (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_write),       //                                         .write
		.Char_Buffer_avalon_char_buffer_slave_read          (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_read),        //                                         .read
		.Char_Buffer_avalon_char_buffer_slave_readdata      (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_readdata),    //                                         .readdata
		.Char_Buffer_avalon_char_buffer_slave_writedata     (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_writedata),   //                                         .writedata
		.Char_Buffer_avalon_char_buffer_slave_byteenable    (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_byteenable),  //                                         .byteenable
		.Char_Buffer_avalon_char_buffer_slave_waitrequest   (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_waitrequest), //                                         .waitrequest
		.Char_Buffer_avalon_char_buffer_slave_chipselect    (mm_interconnect_0_char_buffer_avalon_char_buffer_slave_chipselect),  //                                         .chipselect
		.Char_Buffer_avalon_char_control_slave_address      (mm_interconnect_0_char_buffer_avalon_char_control_slave_address),    //    Char_Buffer_avalon_char_control_slave.address
		.Char_Buffer_avalon_char_control_slave_write        (mm_interconnect_0_char_buffer_avalon_char_control_slave_write),      //                                         .write
		.Char_Buffer_avalon_char_control_slave_read         (mm_interconnect_0_char_buffer_avalon_char_control_slave_read),       //                                         .read
		.Char_Buffer_avalon_char_control_slave_readdata     (mm_interconnect_0_char_buffer_avalon_char_control_slave_readdata),   //                                         .readdata
		.Char_Buffer_avalon_char_control_slave_writedata    (mm_interconnect_0_char_buffer_avalon_char_control_slave_writedata),  //                                         .writedata
		.Char_Buffer_avalon_char_control_slave_byteenable   (mm_interconnect_0_char_buffer_avalon_char_control_slave_byteenable), //                                         .byteenable
		.Char_Buffer_avalon_char_control_slave_chipselect   (mm_interconnect_0_char_buffer_avalon_char_control_slave_chipselect), //                                         .chipselect
		.CPU_debug_mem_slave_address                        (mm_interconnect_0_cpu_debug_mem_slave_address),                      //                      CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write                          (mm_interconnect_0_cpu_debug_mem_slave_write),                        //                                         .write
		.CPU_debug_mem_slave_read                           (mm_interconnect_0_cpu_debug_mem_slave_read),                         //                                         .read
		.CPU_debug_mem_slave_readdata                       (mm_interconnect_0_cpu_debug_mem_slave_readdata),                     //                                         .readdata
		.CPU_debug_mem_slave_writedata                      (mm_interconnect_0_cpu_debug_mem_slave_writedata),                    //                                         .writedata
		.CPU_debug_mem_slave_byteenable                     (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                   //                                         .byteenable
		.CPU_debug_mem_slave_waitrequest                    (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                  //                                         .waitrequest
		.CPU_debug_mem_slave_debugaccess                    (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                  //                                         .debugaccess
		.JTAG_avalon_jtag_slave_address                     (mm_interconnect_0_jtag_avalon_jtag_slave_address),                   //                   JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                       (mm_interconnect_0_jtag_avalon_jtag_slave_write),                     //                                         .write
		.JTAG_avalon_jtag_slave_read                        (mm_interconnect_0_jtag_avalon_jtag_slave_read),                      //                                         .read
		.JTAG_avalon_jtag_slave_readdata                    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                  //                                         .readdata
		.JTAG_avalon_jtag_slave_writedata                   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                 //                                         .writedata
		.JTAG_avalon_jtag_slave_waitrequest                 (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),               //                                         .waitrequest
		.JTAG_avalon_jtag_slave_chipselect                  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                //                                         .chipselect
		.Onchip_Memory_s1_address                           (mm_interconnect_0_onchip_memory_s1_address),                         //                         Onchip_Memory_s1.address
		.Onchip_Memory_s1_write                             (mm_interconnect_0_onchip_memory_s1_write),                           //                                         .write
		.Onchip_Memory_s1_readdata                          (mm_interconnect_0_onchip_memory_s1_readdata),                        //                                         .readdata
		.Onchip_Memory_s1_writedata                         (mm_interconnect_0_onchip_memory_s1_writedata),                       //                                         .writedata
		.Onchip_Memory_s1_byteenable                        (mm_interconnect_0_onchip_memory_s1_byteenable),                      //                                         .byteenable
		.Onchip_Memory_s1_chipselect                        (mm_interconnect_0_onchip_memory_s1_chipselect),                      //                                         .chipselect
		.Onchip_Memory_s1_clken                             (mm_interconnect_0_onchip_memory_s1_clken),                           //                                         .clken
		.Pixel_Buffer_avalon_control_slave_address          (mm_interconnect_0_pixel_buffer_avalon_control_slave_address),        //        Pixel_Buffer_avalon_control_slave.address
		.Pixel_Buffer_avalon_control_slave_write            (mm_interconnect_0_pixel_buffer_avalon_control_slave_write),          //                                         .write
		.Pixel_Buffer_avalon_control_slave_read             (mm_interconnect_0_pixel_buffer_avalon_control_slave_read),           //                                         .read
		.Pixel_Buffer_avalon_control_slave_readdata         (mm_interconnect_0_pixel_buffer_avalon_control_slave_readdata),       //                                         .readdata
		.Pixel_Buffer_avalon_control_slave_writedata        (mm_interconnect_0_pixel_buffer_avalon_control_slave_writedata),      //                                         .writedata
		.Pixel_Buffer_avalon_control_slave_byteenable       (mm_interconnect_0_pixel_buffer_avalon_control_slave_byteenable),     //                                         .byteenable
		.RGB_Resampler_avalon_rgb_slave_read                (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_read),              //           RGB_Resampler_avalon_rgb_slave.read
		.RGB_Resampler_avalon_rgb_slave_readdata            (mm_interconnect_0_rgb_resampler_avalon_rgb_slave_readdata),          //                                         .readdata
		.SDRAM_s1_address                                   (mm_interconnect_0_sdram_s1_address),                                 //                                 SDRAM_s1.address
		.SDRAM_s1_write                                     (mm_interconnect_0_sdram_s1_write),                                   //                                         .write
		.SDRAM_s1_read                                      (mm_interconnect_0_sdram_s1_read),                                    //                                         .read
		.SDRAM_s1_readdata                                  (mm_interconnect_0_sdram_s1_readdata),                                //                                         .readdata
		.SDRAM_s1_writedata                                 (mm_interconnect_0_sdram_s1_writedata),                               //                                         .writedata
		.SDRAM_s1_byteenable                                (mm_interconnect_0_sdram_s1_byteenable),                              //                                         .byteenable
		.SDRAM_s1_readdatavalid                             (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                         .readdatavalid
		.SDRAM_s1_waitrequest                               (mm_interconnect_0_sdram_s1_waitrequest),                             //                                         .waitrequest
		.SDRAM_s1_chipselect                                (mm_interconnect_0_sdram_s1_chipselect),                              //                                         .chipselect
		.timer_s1_address                                   (mm_interconnect_0_timer_s1_address),                                 //                                 timer_s1.address
		.timer_s1_write                                     (mm_interconnect_0_timer_s1_write),                                   //                                         .write
		.timer_s1_readdata                                  (mm_interconnect_0_timer_s1_readdata),                                //                                         .readdata
		.timer_s1_writedata                                 (mm_interconnect_0_timer_s1_writedata),                               //                                         .writedata
		.timer_s1_chipselect                                (mm_interconnect_0_timer_s1_chipselect),                              //                                         .chipselect
		.timer_0_s1_address                                 (mm_interconnect_0_timer_0_s1_address),                               //                               timer_0_s1.address
		.timer_0_s1_write                                   (mm_interconnect_0_timer_0_s1_write),                                 //                                         .write
		.timer_0_s1_readdata                                (mm_interconnect_0_timer_0_s1_readdata),                              //                                         .readdata
		.timer_0_s1_writedata                               (mm_interconnect_0_timer_0_s1_writedata),                             //                                         .writedata
		.timer_0_s1_chipselect                              (mm_interconnect_0_timer_0_s1_chipselect),                            //                                         .chipselect
		.WIFI_Serial_Port_avalon_rs232_slave_address        (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_address),      //      WIFI_Serial_Port_avalon_rs232_slave.address
		.WIFI_Serial_Port_avalon_rs232_slave_write          (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_write),        //                                         .write
		.WIFI_Serial_Port_avalon_rs232_slave_read           (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_read),         //                                         .read
		.WIFI_Serial_Port_avalon_rs232_slave_readdata       (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_readdata),     //                                         .readdata
		.WIFI_Serial_Port_avalon_rs232_slave_writedata      (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_writedata),    //                                         .writedata
		.WIFI_Serial_Port_avalon_rs232_slave_byteenable     (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_byteenable),   //                                         .byteenable
		.WIFI_Serial_Port_avalon_rs232_slave_chipselect     (mm_interconnect_0_wifi_serial_port_avalon_rs232_slave_chipselect)    //                                         .chipselect
	);

	test_irq_mapper irq_mapper (
		.clk           (sys_clk_sys_clk_clk),            //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (sys_clk_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (video_clk_vga_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sys_clk_sys_clk_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.reset_in2      (video_clk_reset_source_reset),       // reset_in2.reset
		.clk            (video_clk_vga_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (sys_clk_reset_source_reset),         // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
